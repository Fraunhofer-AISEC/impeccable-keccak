--Copyright 2024 Fraunhofer Institute for Applied and Integrated Security (AISEC).

--Licensed under the Apache License, Version 2.0 (the "License");
--you may not use this file except in compliance with the License.
--You may obtain a copy of the License at

--    http://www.apache.org/licenses/LICENSE-2.0

--Unless required by applicable law or agreed to in writing, software
--distributed under the License is distributed on an "AS IS" BASIS,
--WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--See the License for the specific language governing permissions and
--limitations under the License.

library work;
	use work.keccak_globals.all;
	use work.keccak_rho_constants.all;

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_arith.all;
	use ieee.std_logic_misc.all;

entity rho_l4 is
	port(
		rho_in : in  k_state;
		rho_out: out k_state
	);
end rho_l4;

--instead of rho_l4_imod4 modules, rho_i matrices can be used, 
--which are stored in keccak_rho_constants.vhd
--that is generated by gen_rho_matrices.py

architecture Behavioural of rho_l4 is
begin
	
	rho_l4_0: for i in 0 to 63 generate
		rho_out(0)(0)(i)<=rho_in(0)(0)(i);
	end generate;
        
	rho_l4_1: for i in 0 to 15 generate
		rho_out(0)(1)(i)<=XOR_REDUCE(rho_in(0)(1) and rho_1(i));
		--m_rho_l4_1mod4 : entity work.rho_l4_1mod4 port map (
		--					data_in => rho_in(0)(1)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(0)(1)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(0)(1)((4*(i+1)-1+4) mod 64 downto (4*i + 4) mod 64)
		--				);
	end generate;
        
	rho_l4_62_01: for i in 0 to 15 generate
		rho_out(0)(2)(i)<=XOR_REDUCE(rho_in(0)(2) and rho_62(i));
		--m_rho_l4_62mod4 : entity work.rho_l4_2mod4 port map (
		--					data_in => rho_in(0)(2)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(0)(2)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(0)(2)((4*(i+1)-1) mod 64 downto (4*i) mod 64)
		--				);
	end generate;
        
	rho_l4_28: for i in 0 to 63 generate
		rho_out(0)(3)(i)<=rho_in(0)(3)((i-28)mod 64);
	end generate;
        
	rho_l4_27: for i in 0 to 15 generate
		rho_out(0)(4)(i)<=XOR_REDUCE(rho_in(0)(4) and rho_27(i));
		--m_rho_l4_27mod4 : entity work.rho_l4_3mod4 port map (
		--					data_in => rho_in(0)(4)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(0)(4)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(0)(4)((4*(i+1)-1+28) mod 64 downto (4*i+28) mod 64)
		--				); 
	end generate;
        
	rho_l4_36: for i in 0 to 63 generate
		rho_out(1)(0)(i)<=rho_in(1)(0)((i-36)mod 64);
	end generate;
        
	rho_44: for i in 0 to 63 generate
		rho_out(1)(1)(i)<=rho_in(1)(1)((i-44)mod 64);
	end generate;
        
	rho_l4_6: for i in 0 to 15 generate
		rho_out(1)(2)(i)<=XOR_REDUCE(rho_in(1)(2) and rho_6(i));
		--m_rho_l4_6mod4 : entity work.rho_l4_2mod4 port map (
		--					data_in => rho_in(1)(2)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(1)(2)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(1)(2)((4*(i+1)-1+8) mod 64 downto (4*i+8) mod 64)
		--				);
	end generate;
        
	rho_l4_55: for i in 0 to 15 generate
		rho_out(1)(3)(i)<=XOR_REDUCE(rho_in(1)(3) and rho_55(i));
		--m_rho_l4_55mod4 : entity work.rho_l4_3mod4 port map (
		--					data_in => rho_in(1)(3)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(1)(3)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(1)(3)((4*(i+1)-1+56) mod 64 downto (4*i+56) mod 64)
		--				); 
	end generate;
        
	rho_l4_20: for i in 0 to 63 generate
		rho_out(1)(4)(i)<=rho_in(1)(4)((i-20)mod 64);
	end generate;

	rho_l4_3: for i in 0 to 15 generate
		rho_out(2)(0)(i)<=XOR_REDUCE(rho_in(2)(0) and rho_3(i));
		--m_rho_l4_3mod4 : entity work.rho_l4_3mod4 port map (
		--					data_in => rho_in(2)(0)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(2)(0)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(2)(0)((4*(i+1)-1+4) mod 64 downto (4*i+4) mod 64)
		--				); 
	end generate;	
        
	rho_l4_10: for i in 0 to 15 generate
		rho_out(2)(1)(i)<=XOR_REDUCE(rho_in(2)(1) and rho_10(i));
		--m_rho_l4_10mod4 : entity work.rho_l4_2mod4 port map (
		--					data_in => rho_in(2)(1)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(2)(1)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(2)(1)((4*(i+1)-1+12) mod 64 downto (4*i+12) mod 64)
		--				);
	end generate;
        
	rho_l4_43: for i in 0 to 15 generate
		rho_out(2)(2)(i)<=XOR_REDUCE(rho_in(2)(2) and rho_43(i));
		--m_rho_l4_43mod4 : entity work.rho_l4_3mod4 port map (
		--					data_in => rho_in(2)(2)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(2)(2)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(2)(2)((4*(i+1)-1+44) mod 64 downto (4*i+44) mod 64)
		--				); 
	end generate;
        
	rho_l4_25: for i in 0 to 15 generate
		rho_out(2)(3)(i)<=XOR_REDUCE(rho_in(2)(3) and rho_25(i));
		--m_rho_l4_25mod4 : entity work.rho_l4_1mod4 port map (
		--					data_in => rho_in(2)(3)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(2)(3)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(2)(3)((4*(i+1)-1+28) mod 64 downto (4*i+28) mod 64)
		--				);
	end generate;
        
	rho_l4_39: for i in 0 to 15 generate
		rho_out(2)(4)(i)<=XOR_REDUCE(rho_in(2)(4) and rho_39(i));
		--m_rho_l4_39mod4 : entity work.rho_l4_3mod4 port map (
		--					data_in => rho_in(2)(4)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(2)(4)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(2)(4)((4*(i+1)-1+40) mod 64 downto (4*i+40) mod 64)
		--				); 
	end generate;
        
	rho_l4_41: for i in 0 to 15 generate
		rho_out(3)(0)(i)<=XOR_REDUCE(rho_in(3)(0) and rho_41(i));
		--m_rho_l4_41mod4 : entity work.rho_l4_1mod4 port map (
		--					data_in => rho_in(3)(0)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(3)(0)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(3)(0)((4*(i+1)-1+44) mod 64 downto (4*i+44) mod 64)
		--				);
	end generate;	
        
	rho_l4_45: for i in 0 to 15 generate
		rho_out(3)(1)(i)<=XOR_REDUCE(rho_in(3)(1) and rho_45(i));
		--m_rho_l4_45mod4 : entity work.rho_l4_1mod4 port map (
		--					data_in => rho_in(3)(1)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(3)(1)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(3)(1)((4*(i+1)-1+48) mod 64 downto (4*i+48) mod 64)
		--				);
	end generate;
        
	rho_l4_15: for i in 0 to 15 generate
		rho_out(3)(2)(i)<=XOR_REDUCE(rho_in(3)(2) and rho_15(i));
		--m_rho_l4_15mod4 : entity work.rho_l4_3mod4 port map (
		--					data_in => rho_in(3)(2)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(3)(2)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(3)(2)((4*(i+1)-1+16) mod 64 downto (4*i+16) mod 64)
		--				); 
	end generate;
        
	rho_l4_21: for i in 0 to 15 generate
		rho_out(3)(3)(i)<=XOR_REDUCE(rho_in(3)(3) and rho_21(i));
		--m_rho_l4_21mod4 : entity work.rho_l4_1mod4 port map (
		--					data_in => rho_in(3)(3)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(3)(3)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(3)(3)((4*(i+1)-1+24) mod 64 downto (4*i+24) mod 64)
		--				);
	end generate;

	rho_l4_8: for i in 0 to 63 generate
		rho_out(3)(4)(i)<=rho_in(3)(4)((i-8)mod 64);
	end generate;

	rho_l4_18: for i in 0 to 15 generate
		rho_out(4)(0)(i)<=XOR_REDUCE(rho_in(4)(0) and rho_18(i));
		--m_rho_l4_18mod4 : entity work.rho_l4_2mod4 port map (
		--					data_in => rho_in(4)(0)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(4)(0)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(4)(0)((4*(i+1)-1+20) mod 64 downto (4*i+20) mod 64)
		--				);
	end generate;	
        
	rho_l4_2: for i in 0 to 15 generate
		rho_out(4)(1)(i)<=XOR_REDUCE(rho_in(4)(1) and rho_2(i));
		--m_rho_l4_2mod4 : entity work.rho_l4_2mod4 port map (
		--					data_in => rho_in(4)(1)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(4)(1)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(4)(1)((4*(i+1)-1+4) mod 64 downto (4*i+4) mod 64)
		--				);
	end generate;
        
	rho_l4_61: for i in 0 to 15 generate
		rho_out(4)(2)(i)<=XOR_REDUCE(rho_in(4)(2) and rho_61(i));
		--m_rho_l4_61mod4 : entity work.rho_l4_1mod4 port map (
		--					data_in => rho_in(4)(2)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(4)(2)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(4)(2)((4*(i+1)-1) mod 64 downto (4*i) mod 64)
		--				);
	end generate;

	rho_l4_56: for i in 0 to 63 generate
		rho_out(4)(3)(i)<=rho_in(4)(3)((i-56)mod 64);
	end generate;
        
	rho_l4_14: for i in 0 to 15 generate
		rho_out(4)(4)(i)<=XOR_REDUCE(rho_in(4)(4) and rho_14(i));
		--m_rho_l4_14mod4 : entity work.rho_l4_2mod4 port map (
		--					data_in => rho_in(4)(4)((4*(i+2)-1) mod 64 downto (4*(i+1)) mod 64) & rho_in(4)(4)(4*(i+1)-1 downto 4*i),
		--					data_out => rho_out(4)(4)((4*(i+1)-1+16) mod 64 downto (4*i+16) mod 64)
		--				);
	end generate;
end Behavioural;
